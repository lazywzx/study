`timescale 1ns / 1ps
module bin_bcd(
clk,rst_n,bin,bcd
    );
	 
input  clk,rst_n;
input  [19:0] bin;
output [23:0] bcd;

reg    [3:0] one,ten,hun,tho,wan,sw;
integer I;
reg    [43:0]shift_reg=44'b0;

////////////////////// 二进制转换为十进制 /////////////////
always @ (posedge clk or negedge rst_n )
begin
shift_reg={23'b0, bin};
	if ( !rst_n )
		  begin
			 one<=0;
			 ten<=0;
			 hun<=0;
			 tho<=0;
			 wan<=0;
			 sw<=0; 
		  end
   else 
	begin 
	   for (I=1; I<=19; I=I+1)
		  begin
				  shift_reg=shift_reg << 1; 
				  
				  if (shift_reg[23:20]+4'b0011>4'b0111)
					  begin
						 shift_reg[23:20]=shift_reg[23:20]+4'b0011; // >7则加3
					  end 
				  if (shift_reg[27:24]+4'b0011>4'b0111)
					  begin
						 shift_reg[27:24]=shift_reg[27:24]+4'b0011;
					  end 
				  if (shift_reg[31:28]+4'b0011>4'b0111)
					  begin
						 shift_reg[31:28]=shift_reg[31:28]+4'b0011;
					  end 
				  if (shift_reg[35:32]+4'b0011>4'b0111)
					  begin
						 shift_reg[35:32]=shift_reg[35:32]+4'b0011;
					  end 
				  if (shift_reg[39:36]+4'b0011>4'b0111)
					  begin
						 shift_reg[39:36]=shift_reg[39:36]+4'b0011;
					  end 
				  if (shift_reg[43:40]+4'b0011>4'b0111)
					  begin
						 shift_reg[43:40]=shift_reg[43:40]+4'b0011;
					  end 		  
				  
		   end
	shift_reg=shift_reg << 1; 
	sw <= shift_reg[43:40];
	wan <= shift_reg[39:36];
	tho <= shift_reg[35:32];
	hun <= shift_reg[31:28];
	ten <= shift_reg[27:24];
	one <= shift_reg[23:20];
	end

end




assign bcd[23:20] = sw;
assign bcd[19:16] = wan;
assign bcd[15:12] = tho;
assign bcd[11:8] = hun;
assign bcd[7:4] = ten;
assign bcd[3:0] = one;

endmodule
